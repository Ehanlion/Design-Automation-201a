/w/home.19/ee/ugrad/palatics/ee201a/lab4/NangateOpenCellLibrary.lef